package my_testbench_pkg;
  import uvm_pkg::*;

  `include "my_transaction.svh"
  `include "my_sequence.svh"
  `include "my_driver.svh"
  `include "my_agent.svh"
  `include "my_env.svh"
  `include "my_test.svh"

endpackage : my_testbench_pkg
